module mem(
    input rst,
    input clk,
    input wire waddr
);

endmodule